-- This file is part of bladeRF-wiphy.
--
-- Copyright (C) 2020 Nuand, LLC.
--
-- This program is free software; you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation; either version 2 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License along
-- with this program; if not, write to the Free Software Foundation, Inc.,
-- 51 Franklin Street, Fifth Floor, Boston, MA 02110-1301 USA.

library ieee ;
    use ieee.std_logic_1164.all ;

library work ;
    use work.wlan_p.all ;

package wlan_tables_p is

    -- Table L-1: MAC PDU Data
    constant TABLE_L_1 : integer_array_t := (
        16#04#, 16#02#, 16#00#, 16#2E#, 16#00#,
        16#60#, 16#08#, 16#CD#, 16#37#, 16#A6#,
        16#00#, 16#20#, 16#D6#, 16#01#, 16#3C#,
        16#F1#, 16#00#, 16#60#, 16#08#, 16#AD#,
        16#3B#, 16#AF#, 16#00#, 16#00#, 16#4A#,
        16#6F#, 16#79#, 16#2C#, 16#20#, 16#62#,
        16#72#, 16#69#, 16#67#, 16#68#, 16#74#,
        16#20#, 16#73#, 16#70#, 16#61#, 16#72#,
        16#6B#, 16#20#, 16#6F#, 16#66#, 16#20#,
        16#64#, 16#69#, 16#76#, 16#69#, 16#6E#,
        16#69#, 16#74#, 16#79#, 16#2C#, 16#0A#,
        16#44#, 16#61#, 16#75#, 16#67#, 16#68#,
        16#74#, 16#65#, 16#72#, 16#20#, 16#6F#,
        16#66#, 16#20#, 16#45#, 16#6C#, 16#79#,
        16#73#, 16#69#, 16#75#, 16#6D#, 16#2C#,
        16#0A#, 16#46#, 16#69#, 16#72#, 16#65#,
        16#2D#, 16#69#, 16#6E#, 16#73#, 16#69#,
        16#72#, 16#65#, 16#64#, 16#20#, 16#77#,
        16#65#, 16#20#, 16#74#, 16#72#, 16#65#,
        16#61#
    ) ;

    -- bladeRF Beacon Frame
    constant BEACON_FRAME : integer_array_t := (
        16#80#, 16#00#, 16#00#, 16#00#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#02#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#,
        16#02#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#dd#, 16#70#, 16#1b#, 16#1e#, 16#78#, 16#01#, 16#05#, 16#00#,
        16#64#, 16#00#, 16#01#, 16#04#, 16#00#, 16#10#, 16#62#, 16#6c#, 16#61#, 16#64#, 16#65#, 16#52#, 16#46#, 16#77#, 16#6c#, 16#61#,
        16#6e#, 16#5f#, 16#53#, 16#53#, 16#49#, 16#44#, 16#01#, 16#08#, 16#82#, 16#84#, 16#8b#, 16#96#, 16#0c#, 16#12#, 16#18#, 16#24#,
        16#03#, 16#01#, 16#01#, 16#05#, 16#04#, 16#01#, 16#02#, 16#00#, 16#00#, 16#2a#, 16#01#, 16#04#, 16#32#, 16#04#, 16#30#, 16#48#,
        16#60#, 16#6c#, 16#7f#, 16#08#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#00#, 16#40#, 16#dd#, 16#18#, 16#00#, 16#50#,
        16#f2#, 16#02#, 16#01#, 16#01#, 16#00#, 16#00#, 16#03#, 16#a4#, 16#00#, 16#00#, 16#27#, 16#a4#, 16#00#, 16#00#, 16#42#, 16#43#,
        16#5e#, 16#00#, 16#62#, 16#32#, 16#2f#, 16#00#, 16#ee#, 16#f7#, 16#d7#, 16#6b#
    ) ;

    constant MIND_FRAME : integer_array_t := (
16#88#, 16#02#, 16#3c#, 16#00#,
16#90#, 16#b6#, 16#86#, 16#e8#,
16#e2#, 16#2f#, 16#00#, 16#1c#,
16#f0#, 16#c5#, 16#e6#, 16#4d#,
16#00#, 16#1c#, 16#f0#, 16#c5#,
16#e6#, 16#4d#, 16#70#, 16#0b#,
16#00#, 16#00#, 16#aa#, 16#aa#,
16#36#, 16#37#
    ) ;

    -- Table L-13: Pre-scrambled data
    constant TABLE_L_13 : integer_array_t := (
        16#00#, 16#00#, 16#04#,
        16#02#, 16#00#, 16#2e#,
        16#00#, 16#60#, 16#08#,
        16#cd#, 16#37#, 16#a6#,
        16#00#, 16#20#, 16#d6#,
        16#01#, 16#3c#, 16#f1#,
        16#00#, 16#60#, 16#08#,
        16#ad#, 16#3b#, 16#af#,
        16#00#, 16#00#, 16#4a#,
        16#6f#, 16#79#, 16#2c#,
        16#20#, 16#62#, 16#72#,
        16#69#, 16#67#, 16#68#,
        16#74#, 16#20#, 16#73#,
        16#70#, 16#61#, 16#72#,
        16#6b#, 16#20#, 16#6f#,
        16#66#, 16#20#, 16#64#,
        16#69#, 16#76#, 16#69#,
        16#6e#, 16#69#, 16#74#,
        16#79#, 16#2c#, 16#0a#,
        16#44#, 16#61#, 16#75#,
        16#67#, 16#68#, 16#74#,
        16#65#, 16#72#, 16#20#,
        16#6f#, 16#66#, 16#20#,
        16#45#, 16#6c#, 16#79#,
        16#73#, 16#69#, 16#75#,
        16#6d#, 16#2c#, 16#0a#,
        16#46#, 16#69#, 16#72#,
        16#65#, 16#2d#, 16#69#,
        16#6e#, 16#73#, 16#69#,
        16#72#, 16#65#, 16#64#,
        16#20#, 16#77#, 16#65#,
        16#20#, 16#74#, 16#72#,
        16#65#, 16#61#, 16#67#,
        16#33#, 16#21#, 16#b6#,
        16#00#, 16#00#, 16#00#,
        16#00#, 16#00#, 16#00#
    ) ;

    -- Post-scrambled data
    constant TABLE_L_15 : integer_array_t := (
        16#6c#, 16#19#, 16#89#,
        16#8f#, 16#68#, 16#21#,
        16#f4#, 16#a5#, 16#61#,
        16#4f#, 16#d7#, 16#ae#,
        16#24#, 16#0c#, 16#f3#,
        16#3a#, 16#e4#, 16#bc#,
        16#53#, 16#98#, 16#c0#,
        16#1e#, 16#35#, 16#b3#,
        16#e3#, 16#f8#, 16#25#,
        16#60#, 16#d6#, 16#25#,
        16#35#, 16#33#, 16#fe#,
        16#f0#, 16#41#, 16#2b#,
        16#8f#, 16#53#, 16#1c#,
        16#83#, 16#41#, 16#be#,
        16#39#, 16#28#, 16#66#,
        16#44#, 16#66#, 16#cd#,
        16#f6#, 16#a3#, 16#d8#,
        16#0d#, 16#d4#, 16#81#,
        16#3b#, 16#2f#, 16#df#,
        16#c3#, 16#58#, 16#f7#,
        16#c6#, 16#52#, 16#eb#,
        16#70#, 16#8f#, 16#9e#,
        16#6a#, 16#90#, 16#81#,
        16#fd#, 16#7c#, 16#a9#,
        16#d1#, 16#55#, 16#12#,
        16#04#, 16#74#, 16#d9#,
        16#e9#, 16#3b#, 16#cd#,
        16#93#, 16#8d#, 16#7b#,
        16#7c#, 16#70#, 16#02#,
        16#20#, 16#99#, 16#a1#,
        16#7d#, 16#8a#, 16#27#,
        16#17#, 16#39#, 16#15#,
        16#a0#, 16#ec#, 16#95#,
        16#16#, 16#91#, 16#10#,
        16#00#, 16#dc#, 16#7f#,
        16#0e#, 16#f2#, 16#c9#
    ) ;

    -- Post Viterbi Encoded (R=3/4) data
    constant TABLE_L_16 : integer_array_t := (
        16#2b#, 16#08#, 16#a1#, 16#f0#,
        16#9d#, 16#b5#, 16#9a#, 16#1d#,
        16#4a#, 16#fb#, 16#e8#, 16#c2#,
        16#8f#, 16#c0#, 16#c8#, 16#73#,
        16#c0#, 16#43#, 16#e0#, 16#19#,
        16#e0#, 16#d3#, 16#eb#, 16#b2#,
        16#af#, 16#98#, 16#fd#, 16#59#,
        16#0f#, 16#8b#, 16#69#, 16#66#,
        16#0c#, 16#aa#, 16#d9#, 16#10#,
        16#56#, 16#8b#, 16#a6#, 16#40#,
        16#64#, 16#b3#, 16#21#, 16#9e#,
        16#8e#, 16#91#, 16#c1#, 16#05#,
        16#b7#, 16#b7#, 16#c5#, 16#d8#,
        16#80#, 16#2f#, 16#a2#, 16#dd#,
        16#6f#, 16#2b#, 16#97#, 16#61#,
        16#d9#, 16#dd#, 16#0d#, 16#12#,
        16#76#, 16#27#, 16#02#, 16#4c#,
        16#92#, 16#bc#, 16#12#, 16#4b#,
        16#6a#, 16#f7#, 16#70#, 16#23#,
        16#27#, 16#8e#, 16#01#, 16#b4#,
        16#d6#, 16#c3#, 16#6a#, 16#60#,
        16#4d#, 16#4b#, 16#cb#, 16#51#,
        16#9c#, 16#b0#, 16#80#, 16#eb#,
        16#89#, 16#34#, 16#14#, 16#40#,
        16#6c#, 16#9e#, 16#2c#, 16#51#,
        16#4b#, 16#7c#, 16#69#, 16#11#,
        16#15#, 16#86#, 16#fd#, 16#be#,
        16#5e#, 16#f9#, 16#be#, 16#28#,
        16#ef#, 16#ca#, 16#55#, 16#03#,
        16#fd#, 16#26#, 16#91#, 16#3b#,
        16#95#, 16#ec#, 16#5b#, 16#23#,
        16#99#, 16#5f#, 16#28#, 16#3e#,
        16#d4#, 16#e9#, 16#f7#, 16#b8#,
        16#13#, 16#75#, 16#8e#, 16#f2#,
        16#a0#, 16#1b#, 16#6c#, 16#e9#,
        16#07#, 16#5d#, 16#b0#, 16#bf#
    ) ;

    -- Table L-19: Data to be modulated
    constant TABLE_L_19 : std_logic_vector(287 downto 0) :=
        x"00000000" &   -- 287 downto 256
        x"00000000" &   -- 255 downto 224
        x"00000000" &   -- 223 downto 192
        x"B6CDB000" &   -- 191 downto 160
        x"C219D6D8" &   -- 159 downto 128
        x"96AF1C76" &   -- 127 downto 96
        x"48B85908" &   -- 95 downto 64
        x"88FD00CE" &   -- 63 downto 32
        x"23F70FEE" ;   -- 32 downto 0

end package ;

